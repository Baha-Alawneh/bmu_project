// BMU UVM Package

package bmu_pkg;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "bmu_seq_item.sv"
  `include "bmu_sequencer.sv"
  `include "bmu_driver.sv"
  `include "bmu_monitor.sv"
  `include "bmu_agent.sv"
  `include "bmu_scoreboard.sv"
  `include "bmu_subscriber.sv"
  `include "bmu_env.sv"
  `include "bmu_base_sequence.sv"
  
  
  `include "sequences/bmu_or_sequence.sv"
  `include "sequences/bmu_orn_sequence.sv"
  `include "sequences/bmu_xor_sequence.sv"
  `include "sequences/bmu_xnor_sequence.sv"
  
  `include "sequences/bmu_srl_sequence.sv"
  `include "sequences/bmu_sra_sequence.sv"
  `include "sequences/bmu_ror_sequence.sv"
  `include "sequences/bmu_binv_sequence.sv"
  `include "sequences/bmu_sh2add_sequence.sv"
  
  `include "sequences/bmu_sub_sequence.sv"
  
  `include "sequences/bmu_sltu_sequence.sv"
  `include "sequences/bmu_slt_sequence.sv"
  `include "sequences/bmu_ctz_sequence.sv"
  `include "sequences/bmu_cpop_sequence.sv"
  `include "sequences/bmu_sext_b_sequence.sv"
  `include "sequences/bmu_max_sequence.sv"
  `include "sequences/bmu_pack_sequence.sv"
  `include "sequences/bmu_grev_sequence.sv"
  
  `include "sequences/bmu_csr_write_sequence.sv"
  `include "sequences/bmu_csr_read_sequence.sv"
  
  `include "sequences/bmu_conflict_sequence.sv"
  
  `include "sequences/bmu_random_sequence.sv"
  
  `include "tests/bmu_base_test.sv"
  `include "tests/bmu_logical_test.sv"
  `include "tests/bmu_shift_test.sv"
  `include "tests/bmu_arithmetic_test.sv"
  `include "tests/bmu_bitmanipulation_test.sv"
  `include "tests/bmu_csr_test.sv"
  `include "tests/bmu_error_test.sv"
  `include "tests/bmu_random_test.sv"
  `include "tests/bmu_regression_test.sv"
  
endpackage : bmu_pkg
